module main

import os { input }

fn main() {
	mut name := input('What is your name: ')
	println('Hello, $name !')
}
